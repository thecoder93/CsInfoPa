** circuit file for profile: simulation 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000us 0 
.OPTIONS DIGINITSTATE= 0
.OPTIONS DIGMNTYMX= 4
.PROBE 
.INC "monostabile-SCHEMATIC1.net" 

.INC "monostabile-SCHEMATIC1.als"


.END
