** circuit file for profile: sim 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000us 0 
.OPTIONS DIGINITSTATE= 0
.PROBE 
.INC "transitionfinder-SCHEMATIC1.net" 

.INC "transitionfinder-SCHEMATIC1.als"


.END
