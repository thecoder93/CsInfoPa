** circuit file for profile: sim 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 160us 0 
.OPTIONS DIGINITSTATE= 0
.PROBE 
.INC "gatedoscillator-SCHEMATIC1.net" 

.INC "gatedoscillator-SCHEMATIC1.als"


.END
