** circuit file for profile: sim 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
.STMLIB ".\PR_ENCODER.stl" 
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500us 0 
.PROBE 
.INC "pr_encoder-SCHEMATIC1.net" 

.INC "pr_encoder-SCHEMATIC1.als"


.END
